`timescale 1ns/1ns
`include "insMem.v"

module insMem_tb;
reg clk;
reg [31:0][0:31]r;
reg l;
reg e;
reg [31:0]address;
wire [31:0][0:0]q;
integer i;


insMem UUT ( .r(r),
 .l(l),
  .address(address),
   .clk(clk),
    .q(q),
    .e(e));

initial begin
    $dumpfile("insMem_tb.vcd");
    $dumpvars(0, insMem_tb);

    // clk= 0;
    // e=0;
    // #10;
    // l = 1;
    // address = 0;
    // r[0] = 32'b00001111000011110000111100001110;
    // r[1] = 32'b00001100000011000000110000001100;
    // for (i = 31; i>1; i--) begin
    //     r[i] = 32'b10000000000000000000000000000000;
    // end
    // clk =1;
    // #10;
    // clk = 0;
    // l=0;
    //     $display("%b", q);
    
    // #10;
    // /////////////////
    // e=1;
    // l = 1;
    // address = 1;
    // r[0] = 32'b00001111000011110000111100001110;
    // r[1] = 32'b00001100000011000000110000001100;
    // for (i = 31; i>1; i--) begin
    //     r[i] = 32'b10000000000000000000000000000000;
    // end
    // clk =1;
    // #10;
    // clk = 0;
    
    //     $display("%b", q);
    
    // #10;
    // //////////////////////////
    // e=0;
    // l = 1;
    // address = 1;
    // r[0] = 32'b00001111000011110000111100001110;
    // r[1] = 32'b00001100000011000000110000001100;
    // for (i = 31; i>1; i--) begin
    //     r[i] = 32'b10000000000000000000000000000000;
    // end
    // clk =1;
    // #10;
    // clk = 0;
    // l=0;
    //     $display("%b", q);
        
    // #10;

    e=1;
    clk=1;
    l=1;
    address = 0;
    r[0] = 32'b00001111000011110000111100001110;
    r[1] = 32'b00001100000011000000110000001100;
    for (i = 30; i>1; i--) begin
        r[i] = 32'b10000000000000000000000000000000;
    end
        r[31] = 32'b11111100000011000000110000001100;
    #10;
    if(q != 32'b00001111000011110000111100001110)
        $display("Error occured in first test");
    ///////////////////

        clk=0;
        l=1;
    #10;
    if(q != 32'b00001111000011110000111100001110)
        $display("Error occured in second test");
    ///////////////////

    clk=1;
    l=1;
    address = 1;
    r[0] = 32'b00001111000011110000111100001110;
    r[1] = 32'b00001100000011000000110000001100;
    for (i = 30; i>1; i--) begin
        r[i] = 32'b10000000000000000000000000000000;
    end
    r[31] = 32'b11111100000011000000110000001100;
    #10;
    if(q != 32'b00001100000011000000110000001100)
        $display("Error occured in third test");
    ///////////////////

        clk=0;
        l=1;
    #10;
    if(q != 32'b00001100000011000000110000001100)
        $display("Error occured in forth test");
    ///////////////////

    clk=1;
    l=0;
    address= 2;
    r[0] = 32'b00001111000011110000111100001110;
    r[1] = 32'b00001100000011000000110000001100;
    for (i = 30; i>1; i--) begin
        r[i] = 32'b10000000000000000000000000000000;
    end
    r[31] = 32'b11111100000011000000110000001100;
    #10;
    if(q != 32'b00001100000011000000110000001100)
        $display("Error occured in fifth test");
    ///////////////////

        clk=0;
        l=0;
    #10;
    if(q != 32'b00001100000011000000110000001100)
        $display("Error occured in sixth test");
    ///////////////////

    clk=1;
    l=1;
    address = 31;
    r[0] = 32'b00001111000011110000111100001110;
    r[1] = 32'b00001100000011000000110000001100;
    for (i = 30; i>1; i--) begin
        r[i] = 32'b10000000000000000000000000000000;
    end
    r[31] = 32'b11111100000011000000110000001100;
    #10;
    if(q != 32'b11111100000011000000110000001100)
        $display("Error occured in seventh test");
    ///////////////////

    clk=0;
    l=1;
    #10;
    if(q != 32'b11111100000011000000110000001100)
        $display("Error occured in eigth test");
    ///////////////////
end

endmodule