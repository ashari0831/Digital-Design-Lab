module insMem ( 
    address, 
    q
);

    reg [31:0][0:31]r;
    input [63:0]address;
    output [31:0][0:0]q;
    integer i;


    initial begin
        r[0] = 32'b00000000111000010010010000100011; //rs2=14, rs1=2, offset[4:0]=8,  SW
        r[4] = 32'b00000000100000010010011100000011;//imm=8, rs1=2, rd=14      LW
        r[8] = 32'b00000000101010011000100100110011;//rs2=10, rs1=19, rd=18       ADD
        r[12] = 32'b01000000101010011000100110110011;// rs2=10, rs1=19, rd=19       SUB
        r[16] = 32'b00000000101010011111101000110011;// rs2=10, rs1=19, rd=20      AND
        r[20] = 32'b00000000101010011110101010110011;// rs2=10, rs1=19, rd=21      OR
        r[24] = 32'b00000000101010011000011101100011;//rs2=10, rs1=19          BEQ
    end
    // initial begin
    //     r[0] = 32'h00000293 ;
    //     r[4] = 32'h00100313 ;
    //     r[8] = 32'h00500393 ;
    //     r[12] =32'h01400E13 ; 
    //     r[16] =32'h0072AEB3 ; 
    //     r[20] =32'h000E8C63 ; 
    //     r[24] =32'h406E0E33 ;
    //     r[28] =  32'h026E0E33;
    //     r[32] = 32'h00128293;
    //     r[36] = 32'hFE5284E3; 
    // end
    
    assign q = r[address];



    
    
endmodule